hola mundo
adoal
module t01pos
enmodule
para comer
necesito pizza
